library verilog;
use verilog.vl_types.all;
entity MPC_GENERATOR_vlg_vec_tst is
end MPC_GENERATOR_vlg_vec_tst;
