library verilog;
use verilog.vl_types.all;
entity ULA_32BIT_vlg_vec_tst is
end ULA_32BIT_vlg_vec_tst;
