library verilog;
use verilog.vl_types.all;
entity MDR_vlg_vec_tst is
end MDR_vlg_vec_tst;
