library verilog;
use verilog.vl_types.all;
entity UNIDADE_CONTROLE_vlg_vec_tst is
end UNIDADE_CONTROLE_vlg_vec_tst;
