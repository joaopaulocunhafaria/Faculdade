library verilog;
use verilog.vl_types.all;
entity decoder2_4_vlg_check_tst is
    port(
        S0              : in     vl_logic;
        S1              : in     vl_logic;
        S2              : in     vl_logic;
        S3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end decoder2_4_vlg_check_tst;
