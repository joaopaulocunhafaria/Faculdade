library verilog;
use verilog.vl_types.all;
entity CONTROL_UNIT_vlg_vec_tst is
end CONTROL_UNIT_vlg_vec_tst;
