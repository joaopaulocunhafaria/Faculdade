library verilog;
use verilog.vl_types.all;
entity REGISTER32bit_vlg_vec_tst is
end REGISTER32bit_vlg_vec_tst;
