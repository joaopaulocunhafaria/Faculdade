library verilog;
use verilog.vl_types.all;
entity OPC_vlg_vec_tst is
end OPC_vlg_vec_tst;
