library verilog;
use verilog.vl_types.all;
entity LV_vlg_vec_tst is
end LV_vlg_vec_tst;
