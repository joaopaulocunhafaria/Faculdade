library verilog;
use verilog.vl_types.all;
entity RAM_TEST_vlg_vec_tst is
end RAM_TEST_vlg_vec_tst;
