library verilog;
use verilog.vl_types.all;
entity MBR_vlg_vec_tst is
end MBR_vlg_vec_tst;
