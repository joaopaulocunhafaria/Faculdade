library verilog;
use verilog.vl_types.all;
entity BANK_REG_vlg_vec_tst is
end BANK_REG_vlg_vec_tst;
