library verilog;
use verilog.vl_types.all;
entity decoder3to8_vlg_vec_tst is
end decoder3to8_vlg_vec_tst;
