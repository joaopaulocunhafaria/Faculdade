library verilog;
use verilog.vl_types.all;
entity REGISTER_4BIT_vlg_vec_tst is
end REGISTER_4BIT_vlg_vec_tst;
