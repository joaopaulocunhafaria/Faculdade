library verilog;
use verilog.vl_types.all;
entity FullAdder_8bit_vlg_vec_tst is
end FullAdder_8bit_vlg_vec_tst;
