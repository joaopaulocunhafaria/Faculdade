library verilog;
use verilog.vl_types.all;
entity H_vlg_vec_tst is
end H_vlg_vec_tst;
