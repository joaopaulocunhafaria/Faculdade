library verilog;
use verilog.vl_types.all;
entity ULA_8bit_vlg_vec_tst is
end ULA_8bit_vlg_vec_tst;
