library verilog;
use verilog.vl_types.all;
entity decoder2to4_vlg_check_tst is
    port(
        s0              : in     vl_logic;
        s1              : in     vl_logic;
        s2              : in     vl_logic;
        s3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end decoder2to4_vlg_check_tst;
