library verilog;
use verilog.vl_types.all;
entity ULA_1BIT_vlg_vec_tst is
end ULA_1BIT_vlg_vec_tst;
