library verilog;
use verilog.vl_types.all;
entity CPP_vlg_vec_tst is
end CPP_vlg_vec_tst;
