library verilog;
use verilog.vl_types.all;
entity TOS_vlg_vec_tst is
end TOS_vlg_vec_tst;
