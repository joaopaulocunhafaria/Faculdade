library verilog;
use verilog.vl_types.all;
entity FullAdder_1bit_vlg_vec_tst is
end FullAdder_1bit_vlg_vec_tst;
