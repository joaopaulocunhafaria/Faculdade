library verilog;
use verilog.vl_types.all;
entity decoder2to4_vlg_vec_tst is
end decoder2to4_vlg_vec_tst;
